** Cascoded common source

.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.param mc_mm_switch=0
.param lx=0.15 wx=162.5 nfx=40 idx=0.5m
.save @m.M1.msky130_fd_pr__nfet_01v8_lvt
.save @m.M2.msky130_fd_pr__nfet_01v8_lvt

* D G S B
M2 out vbias d 0 sky130_fd_pr__nfet_01v8_lvt L={lx} W={wx} nf={nfx} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
M1 d vin 0 0 sky130_fd_pr__nfet_01v8_lvt L={lx} W={wx} nf={nfx} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1

vg  vin  0  0.3
vb  vbias  0  1
is  out  0  {idx}

.control
  op
  *show
  print @m.M1.msky130_fd_pr__nfet_01v8_lvt[gm]
  print @m.M1.msky130_fd_pr__nfet_01v8_lvt[id]
  print @m.M1.msky130_fd_pr__nfet_01v8_lvt[gds]
.endc
.end
